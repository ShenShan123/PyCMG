* instance sweep netlist
X1 d g s e nmos1 L=4e-08 TFIN=2e-08 NFIN=20.0 NRS=1.0 NRD=1.0
.end