* instance sweep netlist
X1 d g s e nmos1 L=2e-08 TFIN=1e-08 NFIN=5.0 NRS=1.0 NRD=1.0
.end