* instance sweep netlist
X1 d g s e nmos1 L=1.6e-08 TFIN=8e-09 NFIN=2.0 NRS=1.0 NRD=1.0
.end