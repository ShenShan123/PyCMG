* Test TSMC7 fixed modelcard syntax
* This test just verifies the file loads and parses correctly

.include "tech_model_cards/TSMC7/cln7_1d8_sp_v1d2_2p2_clean_fixed.l"

* Simple resistor test to verify file loaded
R1 1 0 1k
V1 1 0 1.0

* DC operating point
.op

* End
.end
