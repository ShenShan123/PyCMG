* Test NGSPICE with cleaned TSMC7 modelcard
.include /home/shenshan/pycmg-wrapper/.worktrees/more-techs/build-deep-verify/osdi/bsimcmg.osdi
.lib /home/shenshan/pycmg-wrapper/.worktrees/more-techs/tech_model_cards/TSMC7/cln7_1d8_sp_v1d2_2p2_clean.l Total_svt

* Simple test circuit
* NMOS transistor
M1 drain gate 0 0 nch_svt_mac l=120n nfin=12

* Bias voltages
Vds drain 0 0.5
Vgs gate 0 0.8

* Analysis
.op

* Output
.print dc v(drain) v(gate) i(Vds) i(Vgs)

.end
